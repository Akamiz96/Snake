-------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-------------------------------------------------------------------------------
ENTITY FOOD IS
	PORT	(	clk              :	IN		STD_LOGIC;    
            rst              :	IN		STD_LOGIC
	);
END ENTITY FOOD;
-------------------------------------------------------------------------------
ARCHITECTURE structural OF FOOD IS
	

BEGIN	
	
	

END ARCHITECTURE structural;
------------------------------------------------------------------------------